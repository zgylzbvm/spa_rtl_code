module kos_adder_32 (
    input [31:0] a,b,
    input ci,
    output [31:0] s,
    output co
);

wire [32:0] g[0:5];
wire [31:0] p[0:5];

assign g[0]={a&b,ci};
assign p[0]=a^b;
assign p[1]={p[0][31:31],p[0][30:0]&p[0][31:1]};
assign g[1]={(p[0][31:0]&g[0][31:0])|g[0][32:1],g[0][0:0]};
assign p[2]={p[1][31:29],p[1][28:0]&p[1][30:2]};
assign g[2]={(p[1][30:0]&g[1][30:0])|g[1][32:2],g[1][1:0]};
assign p[3]={p[2][31:25],p[2][24:0]&p[2][28:4]};
assign g[3]={(p[2][28:0]&g[2][28:0])|g[2][32:4],g[2][3:0]};
assign p[4]={p[3][31:17],p[3][16:0]&p[3][24:8]};
assign g[4]={(p[3][24:0]&g[3][24:0])|g[3][32:8],g[3][7:0]};
assign p[5]={p[4][31:1],p[4][0:0]&p[4][16:16]};
assign g[5]={(p[4][16:0]&g[4][16:0])|g[4][32:16],g[4][15:0]};
assign {co,s}={g[5][32]|g[5][0]&p[5][0],p[0]^g[5][31:0]};

endmodule