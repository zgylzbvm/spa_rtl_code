module kos_adder_16 (
    input [15:0] a,b,
    input ci,
    output [15:0] s,
    output co
);

wire [16:0] g[0:4];
wire [15:0] p[0:4];

assign g[0]={a&b,ci};
assign p[0]=a^b;
assign p[1]={p[0][15:15],p[0][14:0]&p[0][15:1]};
assign g[1]={(p[0][15:0]&g[0][15:0])|g[0][16:1],g[0][0:0]};
assign p[2]={p[1][15:13],p[1][12:0]&p[1][14:2]};
assign g[2]={(p[1][14:0]&g[1][14:0])|g[1][16:2],g[1][1:0]};
assign p[3]={p[2][15:9],p[2][8:0]&p[2][12:4]};
assign g[3]={(p[2][12:0]&g[2][12:0])|g[2][16:4],g[2][3:0]};
assign p[4]={p[3][15:1],p[3][0:0]&p[3][8:8]};
assign g[4]={(p[3][8:0]&g[3][8:0])|g[3][16:8],g[3][7:0]};
assign {co,s}={g[4][16]|g[4][0]&p[4][0],p[0]^g[4][15:0]};

endmodule